`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    01:24:19 10/12/2016 
// Design Name: 	Panayiotis Kremmydas
// Module Name:    LEDdecoder 
// Project Name: ???ast???a?? ???as?a 1? - ?d???? ??de???? 7-t�?�?t?? 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module LEDdecoder(input [3:0] char,output [6:0] LED);


//
//G?a t?? ap???d???p???s? t?? 7 s?? 1 t�?�?t?? ???p???ste e?a s??d?ast??? ap???d???p???t?, 
//? ?p???? ?a ??e? ?? e?s?d? t? ??f?? ? ?a?a?t??a p?? ???ete ?a e�fa??sete, ?a? ?a pa???e?
// ?? ???d? t?? t?�?? ?d???s?? t?? 8 t�?�?t??. G?a t?? a?apa??stas? t?? 16 ??f??? apa?te?ta? 
// ?? ???s? a???�?? 4-bit, e?? ta 7 t�?�ata apa?t??? 7 ?e????st? bit (t? de?ad??? ??f??, DP,
// �p??e? ?a �??e? s�?st?, ?d????ta? t? �???�a st? 1).
//
//?ts?, �?a �??f? t?? ap???d???p???t? 7-t�?�?t?? e??a? ? e???:
//
//module LEDdecoder(char, LED);
//input [3:0] char;
//output [6:0] LED;
//
//...
//
//endmodule
//
//S?�p????ste t?? ???p???s? t?? ap???d???p???t? ?a? e????te ?e?t???????, 
//�?s? p??s?�???s??, ?t? ?? t?�?? p?? p????pt??? sta ??f?a t?? LED e??a? ?? 
//?at?????e?, ?a? ????? ?a? t?? s?st? p?????t?ta (0 = a?a��??? ?a? 1 = s�?st?). 
//G?a e?????a st?? epa???e?s?, a??? ?a? ??a t?? ?d???s? t??? st?? p?a??ta, d?a????ste ta ??f?a t?? ap?te??s�at?? 
//LED st?? ?e????st?? e??d??? t?? t�?�?t?? A e?? G.
//
//?ta? ?e???sete ?t? ? ???p???s? e??a? ????, ep?de??te t?? ??d??a Verilog p?? ????ate ?a? ta ap?te??s�ata t?? p??s?�???s?? se ep?t???t? t?? e??ast?????.




endmodule

